LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY n_mem IS
	PORT (
		CS_MEM_IN : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		Rsrc_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		offset_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		ALU_RESULT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RAM_READ_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		PORT_IN_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SP_BUFFERED : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SP_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SP_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		RAM_ADDRESS : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		WB_DATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		RAM_WE : OUT STD_LOGIC
	);
END n_mem;

ARCHITECTURE a_mem OF n_mem IS

	SIGNAL SP_ALU_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PUSH_POP_ADDRESS : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RAM_PORT_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL PushPop_LoadStore : STD_LOGIC;
	SIGNAL SP_AddSubtract : STD_LOGIC;
	SIGNAL MEM_IO : STD_LOGIC;
	SIGNAL PORT_IO : STD_LOGIC;
	SIGNAL READ_WRITE : STD_LOGIC;
BEGIN

	PushPop_LoadStore <= CS_MEM_IN(0);
	SP_AddSubtract <= CS_MEM_IN(1);
	MEM_IO <= CS_MEM_IN(2);
	PORT_IO <= CS_MEM_IN(3);
	READ_WRITE <= CS_MEM_IN(4);

	RAM_WE <= PORT_IO AND READ_WRITE;

	SP_ALU_OUT <= STD_LOGIC_VECTOR(unsigned(SP_IN) + 2) WHEN SP_AddSubtract = '0'
		ELSE
		STD_LOGIC_VECTOR(unsigned(SP_IN) - 2);

	SP_OUT <= SP_ALU_OUT;

	PUSH_POP_ADDRESS <= SP_ALU_OUT WHEN SP_AddSubtract = '0'
		ELSE
		SP_IN;

	RAM_ADDRESS <= PUSH_POP_ADDRESS WHEN PushPop_LoadStore = '0'
		ELSE
		STD_LOGIC_VECTOR(unsigned(Rsrc_IN) + unsigned(offset_IN));

	RAM_PORT_DATA <= PORT_IN_DATA WHEN MEM_IO = '0'
		ELSE
		RAM_READ_DATA;

	WB_DATA <= ALU_RESULT WHEN MEM_IO = '1' OR PORT_IO = '1'
		ELSE
		RAM_PORT_DATA;

END a_mem;