LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY ram IS
GENERIC ( n : integer := 16);
	PORT(
		clk : IN std_logic;
		we  : IN std_logic;
		address : IN  std_logic_vector(2*n-1 DOWNTO 0);
		datain  : IN  std_logic_vector(2*n-1 DOWNTO 0);
		dataout : OUT std_logic_vector(2*n-1 DOWNTO 0));
END ENTITY ram;

ARCHITECTURE syncrama OF ram IS

	TYPE ram_type IS ARRAY(0 TO 2047) OF std_logic_vector(n-1 DOWNTO 0);
	SIGNAL ram : ram_type := (
                0 => "0001000000000001",
		OTHERS => X"0000"
		) ;
	signal RamOut : std_logic_vector(31 DOWNTO 0);
	BEGIN
		PROCESS(clk) IS
			BEGIN
				IF rising_edge(clk) THEN  
					IF we = '1' THEN
						ram(to_integer(unsigned(address))) <= datain;
					END IF;
				END IF;
		END PROCESS;
		RamOut(15 downto 0)<= ram(to_integer(unsigned(address)));
		RamOut(31 downto 16)<= ram(to_integer(unsigned(address))+1);
		dataout <= RamOut;
END syncrama;
